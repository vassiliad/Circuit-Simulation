V1 5 0 2 EXP (2 5 1 0.2 2 0.5)
V2 3 2 0.2
V3 7 6 2
v4 4 8 1 
*SIN (1e-3 0.5 5 1 1 30)
v5 0 6 1 
*PWL(0 1e-3) (1.2 0.1) (1.4 1) (2 0.2) (3 0.4)
r1 1 5 1.5
r2 1 2 1
r3 5 2 50
r4 5 6 0.1
r5 2 6 1.5
r6 3 4 0.1
r7 8 0 1e3
r8 4 0 10

.options  method=be

.tran 0.1 10
.plot V(5) V(1) V(4)
